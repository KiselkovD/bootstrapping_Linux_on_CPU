module test;
    initial $display("hello");
endmodule
